/* AND2 */

module AND2 ( A, B, X );

input wire A, B;
output wire X;

    assign X = A;

endmodule