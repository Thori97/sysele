`define fs 2048
`define N 128
`define logN 7